LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY P_tb1 IS END ENTITY;
ARCHITECTURE ARCH_P_tb1 OF P_tb1 IS
COMPONENT P1 IS PORT (
A :IN STD_LOGIC_VECTOR(7 DOWNTO 0);
Y :OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;
SIGNAL CLK :STD_LOGIC := '0';
SIGNAL A :STD_LOGIC_VECTOR(7 DOWNTO 0) := B"00000000";
SIGNAL Y :STD_LOGIC_VECTOR(7 DOWNTO 0) := B"00000000";
SIGNAL CLKp :time := 40 ns;

BEGIN
uut: permutation PORT MAP (A, Y);
PROCESS
BEGIN
CLK <= '0'; wait for CLKp/2;
CLK <= '1'; wait for CLKp/2;
END PROCESS;
PROCESS
BEGIN
A <= B"00000000"; wait for CLKp;
A <= B"00000001"; wait for CLKp;
A <= B"00000010"; wait for CLKp;
A <= B"00000100"; wait for CLKp;
A <= B"00001000"; wait for CLKp;
A <= B"00010000"; wait for CLKp;
A <= B"00100000"; wait for CLKp;
A <= B"01000000"; wait for CLKp;
A <= B"10000000"; wait for CLKp;
END PROCESS;
END ARCHITECTURE;
mgr