LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY sbox IS PORT
(
DATA_IN :IN STD_LOGIC_VECTOR(47 DOWNTO 0);
DATA_OUT :OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END sbox;
ARCHITECTURE ARCH_sbox OF sbox IS

--type INT_ARRAY is array (31 downto 0) of integer range 0 to 15;
--signal sbox_1 : INT_ARRAY :=(14,4,13,1,2,15,11,8,3,10,6,12,5,9,0,7,0,15,7,4,14,2,13,1,10,6,12,11,9,5,3,8,4,1,14,8,13,6,2,11,15,12,9,7,3,10,5,0,15,12,8,2,4,9,1,7,5,11,3,14,10,0,6,13);
--signal sbox_2 : INT_ARRAY :=(15,1,8,14,6,11,3,4,9,7,2,13,12,0,5,10,3,13,4,7,15,2,8,14,12,0,1,10,6,9,11,5,0,14,7,11,10,4,13,1,5,8,12,6,9,3,2,15,13,8,10,1,3,15,4,2,11,6,7,12,0,5,14,9);
--signal sbox_3 : INT_ARRAY :=(10,0,9,14,6,3,15,5,1,13,12,7,11,4,2,8,13,7,0,9,3,4,6,10,2,8,5,14,12,11,15,1,13,6,4,9,8,15,3,0,11,1,2,12,5,10,14,7,1,10,13,0,6,9,8,7,4,15,14,3,11,5,2,12);
--signal sbox_4 : INT_ARRAY :=(7,13,14,3,0,6,9,10,1,2,8,5,11,12,4,15,13,8,11,5,6,15,0,3,4,7,2,12,1,10,14,9,10,6,9,0,12,11,7,13,15,1,3,14,5,2,8,4,3,15,0,6,10,1,13,8,9,4,5,11,12,7,2,14);
--signal sbox_5 : INT_ARRAY :=(2,12,4,1,7,10,11,6,8,5,3,15,13,0,14,9,14,11,2,12,4,7,13,1,5,0,15,10,3,9,8,6,4,2,1,11,10,13,7,8,15,9,12,5,6,3,0,14,11,8,12,7,1,14,2,13,6,15,0,9,10,4,5,3);
--signal sbox_6 : INT_ARRAY :=(12,1,10,15,9,2,6,8,0,13,3,4,14,7,5,11,10,15,4,2,7,12,9,5,6,1,13,14,0,11,3,8,9,14,15,5,2,8,12,3,7,0,4,10,1,13,11,6,4,3,2,12,9,5,15,10,11,14,1,7,6,0,8,13);
--signal sbox_7 : INT_ARRAY :=(4,11,2,14,15,0,8,13,3,12,9,7,5,10,6,1,13,0,11,7,4,9,1,10,14,3,5,12,2,15,8,6,1,4,11,13,12,3,7,14,10,15,6,8,0,5,9,2,6,11,13,8,1,4,10,7,9,5,0,15,14,2,3,12);
--signal sbox_8 : INT_ARRAY :=(13,2,8,4,6,15,11,1,10,9,3,14,5,0,12,7,1,15,13,8,10,3,7,4,12,5,6,11,0,14,9,2,7,11,4,1,9,12,14,2,0,6,10,13,15,3,5,8,2,1,14,7,4,10,8,13,15,12,9,0,3,5,6,11);

BEGIN
--pierwsze 6 bitów
DATA_OUT(31 downto 28)<=b"1110" when DATA_IN(47 downto 42)=b"000000" else
								b"0000" when DATA_IN(47 downto 42)=b"000001" else
								b"0100" when DATA_IN(47 downto 42)=b"000010" else
								b"1111" when DATA_IN(47 downto 42)=b"000011" else
								b"1101" when DATA_IN(47 downto 42)=b"000100" else
								b"0111" when DATA_IN(47 downto 42)=b"000101" else
								b"0001" when DATA_IN(47 downto 42)=b"000110" else
								b"0100" when DATA_IN(47 downto 42)=b"000111" else
								b"0010" when DATA_IN(47 downto 42)=b"001000" else
								b"1110" when DATA_IN(47 downto 42)=b"001001" else
								b"1111" when DATA_IN(47 downto 42)=b"001010" else
								b"0010" when DATA_IN(47 downto 42)=b"001011" else
								b"1011" when DATA_IN(47 downto 42)=b"001100" else
								b"1101" when DATA_IN(47 downto 42)=b"001101" else
								b"1000" when DATA_IN(47 downto 42)=b"001110" else
								b"0001" when DATA_IN(47 downto 42)=b"001111" else
								b"0011" when DATA_IN(47 downto 42)=b"010000" else
								b"1010" when DATA_IN(47 downto 42)=b"010001" else
								b"1010" when DATA_IN(47 downto 42)=b"010010" else
								b"0110" when DATA_IN(47 downto 42)=b"010011" else
								b"0110" when DATA_IN(47 downto 42)=b"010100" else
								b"1100" when DATA_IN(47 downto 42)=b"010101" else
								b"1100" when DATA_IN(47 downto 42)=b"010110" else
								b"1011" when DATA_IN(47 downto 42)=b"010111" else
								b"0101" when DATA_IN(47 downto 42)=b"011000" else
								b"1001" when DATA_IN(47 downto 42)=b"011001" else
								b"1001" when DATA_IN(47 downto 42)=b"011010" else
								b"0101" when DATA_IN(47 downto 42)=b"011011" else
								b"0000" when DATA_IN(47 downto 42)=b"011100" else
								b"0011" when DATA_IN(47 downto 42)=b"011101" else
								b"0111" when DATA_IN(47 downto 42)=b"011110" else
								b"1000" when DATA_IN(47 downto 42)=b"011111" else
								b"0100" when DATA_IN(47 downto 42)=b"100000" else
								b"1111" when DATA_IN(47 downto 42)=b"100001" else
								b"0001" when DATA_IN(47 downto 42)=b"100010" else
								b"1100" when DATA_IN(47 downto 42)=b"100011" else
								b"1110" when DATA_IN(47 downto 42)=b"100100" else
								b"1000" when DATA_IN(47 downto 42)=b"100101" else
								b"1000" when DATA_IN(47 downto 42)=b"100110" else
								b"0010" when DATA_IN(47 downto 42)=b"100111" else
								b"1101" when DATA_IN(47 downto 42)=b"101000" else
								b"0100" when DATA_IN(47 downto 42)=b"101001" else
								b"0110" when DATA_IN(47 downto 42)=b"101010" else
								b"1001" when DATA_IN(47 downto 42)=b"101011" else
								b"0010" when DATA_IN(47 downto 42)=b"101100" else
								b"0001" when DATA_IN(47 downto 42)=b"101101" else
								b"1011" when DATA_IN(47 downto 42)=b"101110" else
								b"0111" when DATA_IN(47 downto 42)=b"101111" else
								b"1111" when DATA_IN(47 downto 42)=b"110000" else
								b"0101" when DATA_IN(47 downto 42)=b"110001" else
								b"1100" when DATA_IN(47 downto 42)=b"110010" else
								b"1011" when DATA_IN(47 downto 42)=b"110011" else
								b"1001" when DATA_IN(47 downto 42)=b"110100" else
								b"0011" when DATA_IN(47 downto 42)=b"110101" else
								b"0111" when DATA_IN(47 downto 42)=b"110110" else
								b"1110" when DATA_IN(47 downto 42)=b"110111" else
								b"0011" when DATA_IN(47 downto 42)=b"111000" else
								b"1010" when DATA_IN(47 downto 42)=b"111001" else
								b"1010" when DATA_IN(47 downto 42)=b"111010" else
								b"0000" when DATA_IN(47 downto 42)=b"111011" else
								b"0101" when DATA_IN(47 downto 42)=b"111100" else
								b"0110" when DATA_IN(47 downto 42)=b"111101" else
								b"0000" when DATA_IN(47 downto 42)=b"111110" else
								b"1101" when DATA_IN(47 downto 42)=b"111111" else
								(others=>'0');
--drugie 6 bitów
DATA_OUT(27 downto 24)<=B"1111" when DATA_IN(41 downto 36)=b"000000" else
								B"0001" when DATA_IN(41 downto 36)=b"000010" else
								b"1000" when DATA_IN(41 downto 36)=b"000100" else
								b"1110" when DATA_IN(41 downto 36)=b"000110" else
								b"0110" when DATA_IN(41 downto 36)=b"001000" else
								b"1011" when DATA_IN(41 downto 36)=b"001010" else
								b"0011" when DATA_IN(41 downto 36)=b"001100" else
								b"0100" when DATA_IN(41 downto 36)=b"001110" else
								b"1001" when DATA_IN(41 downto 36)=b"010000" else
								b"0111" when DATA_IN(41 downto 36)=b"010010" else
								b"0010" when DATA_IN(41 downto 36)=b"010100" else
								b"1101" when DATA_IN(41 downto 36)=b"010110" else
								b"1100" when DATA_IN(41 downto 36)=b"011000" else
								b"0000" when DATA_IN(41 downto 36)=b"011010" else
								b"0101" when DATA_IN(41 downto 36)=b"011100" else
								b"1010" when DATA_IN(41 downto 36)=b"011110" else
								b"0011" when DATA_IN(41 downto 36)=b"000001" else
								b"1101" when DATA_IN(41 downto 36)=b"000011" else
								b"0100" when DATA_IN(41 downto 36)=b"000101" else
								b"0111" when DATA_IN(41 downto 36)=b"000111" else
								b"1111" when DATA_IN(41 downto 36)=b"001001" else
								b"0010" when DATA_IN(41 downto 36)=b"001011" else
								b"1000" when DATA_IN(41 downto 36)=b"001101" else
								b"1110" when DATA_IN(41 downto 36)=b"001111" else
								b"1100" when DATA_IN(41 downto 36)=b"010001" else
								b"0000" when DATA_IN(41 downto 36)=b"010011" else
								b"0001" when DATA_IN(41 downto 36)=b"010101" else
								b"1010" when DATA_IN(41 downto 36)=b"010111" else
								b"0110" when DATA_IN(41 downto 36)=b"011001" else
								b"1001" when DATA_IN(41 downto 36)=b"011011" else
								b"1011" when DATA_IN(41 downto 36)=b"011101" else
								b"0101" when DATA_IN(41 downto 36)=b"011111" else
								b"0000" when DATA_IN(41 downto 36)=b"100000" else
								b"1110" when DATA_IN(41 downto 36)=b"100010" else
								b"0111" when DATA_IN(41 downto 36)=b"100100" else
								b"1011" when DATA_IN(41 downto 36)=b"100110" else
								b"1010" when DATA_IN(41 downto 36)=b"101000" else
								b"0100" when DATA_IN(41 downto 36)=b"101010" else
								b"1101" when DATA_IN(41 downto 36)=b"101100" else
								b"0001" when DATA_IN(41 downto 36)=b"101110" else
								b"0101" when DATA_IN(41 downto 36)=b"110000" else
								b"1000" when DATA_IN(41 downto 36)=b"110010" else
								b"1100" when DATA_IN(41 downto 36)=b"110100" else
								b"0110" when DATA_IN(41 downto 36)=b"110110" else
								b"1001" when DATA_IN(41 downto 36)=b"111000" else
								b"0011" when DATA_IN(41 downto 36)=b"111010" else
								b"0010" when DATA_IN(41 downto 36)=b"111100" else
								b"1111" when DATA_IN(41 downto 36)=b"111110" else
								b"1101" when DATA_IN(41 downto 36)=b"100001" else
								b"1000" when DATA_IN(41 downto 36)=b"100011" else
								b"1010" when DATA_IN(41 downto 36)=b"100101" else
								b"0001" when DATA_IN(41 downto 36)=b"100111" else
								b"0011" when DATA_IN(41 downto 36)=b"101001" else
								b"1111" when DATA_IN(41 downto 36)=b"101011" else
								b"0100" when DATA_IN(41 downto 36)=b"101101" else
								b"0010" when DATA_IN(41 downto 36)=b"101111" else
								b"1011" when DATA_IN(41 downto 36)=b"110001" else
								b"0110" when DATA_IN(41 downto 36)=b"110011" else
								b"0111" when DATA_IN(41 downto 36)=b"110101" else
								b"1100" when DATA_IN(41 downto 36)=b"110111" else
								b"0000" when DATA_IN(41 downto 36)=b"111001" else
								b"0101" when DATA_IN(41 downto 36)=b"111011" else
								b"1110" when DATA_IN(41 downto 36)=b"111101" else
								b"1001" when DATA_IN(41 downto 36)=b"111111" else
								(others=>'0');
--trzeci sbox		
DATA_OUT(23 downto 20)<=b"1010" when DATA_IN(35 downto 30)=b"000000" else
								b"0000" when DATA_IN(35 downto 30)=b"000010" else
								b"1001" when DATA_IN(35 downto 30)=b"000100" else
								b"1110" when DATA_IN(35 downto 30)=b"000110" else
								b"0110" when DATA_IN(35 downto 30)=b"001000" else
								b"0011" when DATA_IN(35 downto 30)=b"001010" else
								b"1111" when DATA_IN(35 downto 30)=b"001100" else
								b"0101" when DATA_IN(35 downto 30)=b"001110" else
								b"0001" when DATA_IN(35 downto 30)=b"010000" else
								b"1101" when DATA_IN(35 downto 30)=b"010010" else
								b"1100" when DATA_IN(35 downto 30)=b"010100" else
								b"0111" when DATA_IN(35 downto 30)=b"010110" else
								b"1011" when DATA_IN(35 downto 30)=b"011000" else
								b"0100" when DATA_IN(35 downto 30)=b"011010" else
								b"0010" when DATA_IN(35 downto 30)=b"011100" else
								b"1000" when DATA_IN(35 downto 30)=b"011110" else
								b"1101" when DATA_IN(35 downto 30)=b"000001" else
								b"0111" when DATA_IN(35 downto 30)=b"000011" else
								b"0000" when DATA_IN(35 downto 30)=b"000101" else
								b"1001" when DATA_IN(35 downto 30)=b"000111" else
								b"0011" when DATA_IN(35 downto 30)=b"001001" else
								b"0100" when DATA_IN(35 downto 30)=b"001011" else
								b"0110" when DATA_IN(35 downto 30)=b"001101" else
								b"1010" when DATA_IN(35 downto 30)=b"001111" else
								b"0010" when DATA_IN(35 downto 30)=b"010001" else
								b"1000" when DATA_IN(35 downto 30)=b"010011" else
								b"0101" when DATA_IN(35 downto 30)=b"010101" else
								b"1110" when DATA_IN(35 downto 30)=b"010111" else
								b"1100" when DATA_IN(35 downto 30)=b"011001" else
								b"1011" when DATA_IN(35 downto 30)=b"011011" else
								b"1111" when DATA_IN(35 downto 30)=b"011101" else
								b"0001" when DATA_IN(35 downto 30)=b"011111" else
								b"1101" when DATA_IN(35 downto 30)=b"100000" else
								b"0110" when DATA_IN(35 downto 30)=b"100010" else
								b"0100" when DATA_IN(35 downto 30)=b"100100" else
								b"1001" when DATA_IN(35 downto 30)=b"100110" else
								b"1000" when DATA_IN(35 downto 30)=b"101000" else
								b"1111" when DATA_IN(35 downto 30)=b"101010" else
								b"0011" when DATA_IN(35 downto 30)=b"101100" else
								b"0000" when DATA_IN(35 downto 30)=b"101110" else
								b"1011" when DATA_IN(35 downto 30)=b"110000" else
								b"0001" when DATA_IN(35 downto 30)=b"110010" else
								b"0010" when DATA_IN(35 downto 30)=b"110100" else
								b"1100" when DATA_IN(35 downto 30)=b"110110" else
								b"0101" when DATA_IN(35 downto 30)=b"111000" else
								b"1010" when DATA_IN(35 downto 30)=b"111010" else
								b"1110" when DATA_IN(35 downto 30)=b"111100" else
								b"0111" when DATA_IN(35 downto 30)=b"111110" else
								b"0001" when DATA_IN(35 downto 30)=b"100001" else
								b"1010" when DATA_IN(35 downto 30)=b"100011" else
								b"1101" when DATA_IN(35 downto 30)=b"100101" else
								b"0000" when DATA_IN(35 downto 30)=b"100111" else
								b"0110" when DATA_IN(35 downto 30)=b"101001" else
								b"1001" when DATA_IN(35 downto 30)=b"101011" else
								b"1000" when DATA_IN(35 downto 30)=b"101101" else
								b"0111" when DATA_IN(35 downto 30)=b"101111" else
								b"0100" when DATA_IN(35 downto 30)=b"110001" else
								b"1111" when DATA_IN(35 downto 30)=b"110011" else
								b"1110" when DATA_IN(35 downto 30)=b"110101" else
								b"0011" when DATA_IN(35 downto 30)=b"110111" else
								b"1011" when DATA_IN(35 downto 30)=b"111001" else
								b"0101" when DATA_IN(35 downto 30)=b"111011" else
								b"0010" when DATA_IN(35 downto 30)=b"111101" else
								b"1100" when DATA_IN(35 downto 30)=b"111111" else
								(others=>'0');
-- czwarty sbox
DATA_OUT(19 downto 16)<=b"0111" when DATA_IN(29 downto 24)=b"000000" else
								b"1101" when DATA_IN(29 downto 24)=b"000010" else
								b"1110" when DATA_IN(29 downto 24)=b"000100" else
								b"0011" when DATA_IN(29 downto 24)=b"000110" else
								b"0000" when DATA_IN(29 downto 24)=b"001000" else
								b"0110" when DATA_IN(29 downto 24)=b"001010" else
								b"1001" when DATA_IN(29 downto 24)=b"001100" else
								b"1010" when DATA_IN(29 downto 24)=b"001110" else
								b"0001" when DATA_IN(29 downto 24)=b"010000" else
								b"0010" when DATA_IN(29 downto 24)=b"010010" else
								b"1000" when DATA_IN(29 downto 24)=b"010100" else
								b"0101" when DATA_IN(29 downto 24)=b"010110" else
								b"1011" when DATA_IN(29 downto 24)=b"011000" else
								b"1100" when DATA_IN(29 downto 24)=b"011010" else
								b"0100" when DATA_IN(29 downto 24)=b"011100" else
								b"1111" when DATA_IN(29 downto 24)=b"011110" else
								b"1101" when DATA_IN(29 downto 24)=b"000001" else
								b"1000" when DATA_IN(29 downto 24)=b"000011" else
								b"1011" when DATA_IN(29 downto 24)=b"000101" else
								b"0101" when DATA_IN(29 downto 24)=b"000111" else
								b"0110" when DATA_IN(29 downto 24)=b"001001" else
								b"1111" when DATA_IN(29 downto 24)=b"001011" else
								b"0000" when DATA_IN(29 downto 24)=b"001101" else
								b"0011" when DATA_IN(29 downto 24)=b"001111" else
								b"0100" when DATA_IN(29 downto 24)=b"010001" else
								b"0111" when DATA_IN(29 downto 24)=b"010011" else
								b"0010" when DATA_IN(29 downto 24)=b"010101" else
								b"1100" when DATA_IN(29 downto 24)=b"010111" else
								b"0001" when DATA_IN(29 downto 24)=b"011001" else
								b"1010" when DATA_IN(29 downto 24)=b"011011" else
								b"1110" when DATA_IN(29 downto 24)=b"011101" else
								b"1001" when DATA_IN(29 downto 24)=b"011111" else
								b"1010" when DATA_IN(29 downto 24)=b"100000" else
								b"0110" when DATA_IN(29 downto 24)=b"100010" else
								b"1001" when DATA_IN(29 downto 24)=b"100100" else
								b"0000" when DATA_IN(29 downto 24)=b"100110" else
								b"1100" when DATA_IN(29 downto 24)=b"101000" else
								b"1011" when DATA_IN(29 downto 24)=b"101010" else
								b"0111" when DATA_IN(29 downto 24)=b"101100" else
								b"1101" when DATA_IN(29 downto 24)=b"101110" else
								b"1111" when DATA_IN(29 downto 24)=b"110000" else
								b"0001" when DATA_IN(29 downto 24)=b"110010" else
								b"0011" when DATA_IN(29 downto 24)=b"110100" else
								b"1110" when DATA_IN(29 downto 24)=b"110110" else
								b"0101" when DATA_IN(29 downto 24)=b"111000" else
								b"0010" when DATA_IN(29 downto 24)=b"111010" else
								b"1000" when DATA_IN(29 downto 24)=b"111100" else
								b"0100" when DATA_IN(29 downto 24)=b"111110" else
								b"0011" when DATA_IN(29 downto 24)=b"100001" else
								b"1111" when DATA_IN(29 downto 24)=b"100011" else
								b"0000" when DATA_IN(29 downto 24)=b"100101" else
								b"0110" when DATA_IN(29 downto 24)=b"100111" else
								b"1010" when DATA_IN(29 downto 24)=b"101001" else
								b"0001" when DATA_IN(29 downto 24)=b"101011" else
								b"1101" when DATA_IN(29 downto 24)=b"101101" else
								b"1000" when DATA_IN(29 downto 24)=b"101111" else
								b"1001" when DATA_IN(29 downto 24)=b"110001" else
								b"0100" when DATA_IN(29 downto 24)=b"110011" else
								b"0101" when DATA_IN(29 downto 24)=b"110101" else
								b"1011" when DATA_IN(29 downto 24)=b"110111" else
								b"1100" when DATA_IN(29 downto 24)=b"111001" else
								b"0111" when DATA_IN(29 downto 24)=b"111011" else
								b"0010" when DATA_IN(29 downto 24)=b"111101" else
								b"1110" when DATA_IN(29 downto 24)=b"111111" else
								(others=>'0');
--piąty sbox			
DATA_OUT(15 downto 12)<=b"0010" when DATA_IN(23 downto 18)=b"000000" else
								b"1100" when DATA_IN(23 downto 18)=b"000010" else
								b"0100" when DATA_IN(23 downto 18)=b"000100" else
								b"0001" when DATA_IN(23 downto 18)=b"000110" else
								b"0111" when DATA_IN(23 downto 18)=b"001000" else
								b"1010" when DATA_IN(23 downto 18)=b"001010" else
								b"1011" when DATA_IN(23 downto 18)=b"001100" else
								b"0110" when DATA_IN(23 downto 18)=b"001110" else
								b"1000" when DATA_IN(23 downto 18)=b"010000" else
								b"0101" when DATA_IN(23 downto 18)=b"010010" else
								b"0011" when DATA_IN(23 downto 18)=b"010100" else
								b"1111" when DATA_IN(23 downto 18)=b"010110" else
								b"1101" when DATA_IN(23 downto 18)=b"011000" else
								b"0000" when DATA_IN(23 downto 18)=b"011010" else
								b"1110" when DATA_IN(23 downto 18)=b"011100" else
								b"1001" when DATA_IN(23 downto 18)=b"011110" else
								b"1110" when DATA_IN(23 downto 18)=b"000001" else
								b"1011" when DATA_IN(23 downto 18)=b"000011" else
								b"0010" when DATA_IN(23 downto 18)=b"000101" else
								b"1100" when DATA_IN(23 downto 18)=b"000111" else
								b"0100" when DATA_IN(23 downto 18)=b"001001" else
								b"0111" when DATA_IN(23 downto 18)=b"001011" else
								b"1101" when DATA_IN(23 downto 18)=b"001101" else
								b"0001" when DATA_IN(23 downto 18)=b"001111" else
								b"0101" when DATA_IN(23 downto 18)=b"010001" else
								b"0000" when DATA_IN(23 downto 18)=b"010011" else
								b"1111" when DATA_IN(23 downto 18)=b"010101" else
								b"1010" when DATA_IN(23 downto 18)=b"010111" else
								b"0011" when DATA_IN(23 downto 18)=b"011001" else
								b"1001" when DATA_IN(23 downto 18)=b"011011" else
								b"1000" when DATA_IN(23 downto 18)=b"011101" else
								b"0110" when DATA_IN(23 downto 18)=b"011111" else
								b"0100" when DATA_IN(23 downto 18)=b"100000" else
								b"0010" when DATA_IN(23 downto 18)=b"100010" else
								b"0001" when DATA_IN(23 downto 18)=b"100100" else
								b"1011" when DATA_IN(23 downto 18)=b"100110" else
								b"1010" when DATA_IN(23 downto 18)=b"101000" else
								b"1101" when DATA_IN(23 downto 18)=b"101010" else
								b"0111" when DATA_IN(23 downto 18)=b"101100" else
								b"1000" when DATA_IN(23 downto 18)=b"101110" else
								b"1111" when DATA_IN(23 downto 18)=b"110000" else
								b"1001" when DATA_IN(23 downto 18)=b"110010" else
								b"1100" when DATA_IN(23 downto 18)=b"110100" else
								b"0101" when DATA_IN(23 downto 18)=b"110110" else
								b"0110" when DATA_IN(23 downto 18)=b"111000" else
								b"0011" when DATA_IN(23 downto 18)=b"111010" else
								b"0000" when DATA_IN(23 downto 18)=b"111100" else
								b"1110" when DATA_IN(23 downto 18)=b"111110" else
								b"1011" when DATA_IN(23 downto 18)=b"100001" else
								b"1000" when DATA_IN(23 downto 18)=b"100011" else
								b"1100" when DATA_IN(23 downto 18)=b"100101" else
								b"0111" when DATA_IN(23 downto 18)=b"100111" else
								b"0001" when DATA_IN(23 downto 18)=b"101001" else
								b"1110" when DATA_IN(23 downto 18)=b"101011" else
								b"0010" when DATA_IN(23 downto 18)=b"101101" else
								b"1101" when DATA_IN(23 downto 18)=b"101111" else
								b"0110" when DATA_IN(23 downto 18)=b"110001" else
								b"1111" when DATA_IN(23 downto 18)=b"110011" else
								b"0000" when DATA_IN(23 downto 18)=b"110101" else
								b"1001" when DATA_IN(23 downto 18)=b"110111" else
								b"1010" when DATA_IN(23 downto 18)=b"111001" else
								b"0100" when DATA_IN(23 downto 18)=b"111011" else
								b"0101" when DATA_IN(23 downto 18)=b"111101" else
								b"0011" when DATA_IN(23 downto 18)=b"111111" else
								(others=>'0');
--szósty sbox			
DATA_OUT(11 downto 8)<= b"1100" when DATA_IN(17 downto 12)=b"000000" else
								b"0001" when DATA_IN(17 downto 12)=b"000010" else
								b"1010" when DATA_IN(17 downto 12)=b"000100" else
								b"1111" when DATA_IN(17 downto 12)=b"000110" else
								b"1001" when DATA_IN(17 downto 12)=b"001000" else
								b"0010" when DATA_IN(17 downto 12)=b"001010" else
								b"0110" when DATA_IN(17 downto 12)=b"001100" else
								b"1000" when DATA_IN(17 downto 12)=b"001110" else
								b"0000" when DATA_IN(17 downto 12)=b"010000" else
								b"1101" when DATA_IN(17 downto 12)=b"010010" else
								b"0011" when DATA_IN(17 downto 12)=b"010100" else
								b"0100" when DATA_IN(17 downto 12)=b"010110" else
								b"1110" when DATA_IN(17 downto 12)=b"011000" else
								b"0111" when DATA_IN(17 downto 12)=b"011010" else
								b"0101" when DATA_IN(17 downto 12)=b"011100" else
								b"1011" when DATA_IN(17 downto 12)=b"011110" else
								b"1010" when DATA_IN(17 downto 12)=b"000001" else
								b"1111" when DATA_IN(17 downto 12)=b"000011" else
								b"0100" when DATA_IN(17 downto 12)=b"000101" else
								b"0010" when DATA_IN(17 downto 12)=b"000111" else
								b"0111" when DATA_IN(17 downto 12)=b"001001" else
								b"1100" when DATA_IN(17 downto 12)=b"001011" else
								b"1001" when DATA_IN(17 downto 12)=b"001101" else
								b"0101" when DATA_IN(17 downto 12)=b"001111" else
								b"0110" when DATA_IN(17 downto 12)=b"010001" else
								b"0001" when DATA_IN(17 downto 12)=b"010011" else
								b"1101" when DATA_IN(17 downto 12)=b"010101" else
								b"1110" when DATA_IN(17 downto 12)=b"010111" else
								b"0000" when DATA_IN(17 downto 12)=b"011001" else
								b"1011" when DATA_IN(17 downto 12)=b"011011" else
								b"0011" when DATA_IN(17 downto 12)=b"011101" else
								b"1000" when DATA_IN(17 downto 12)=b"011111" else
								b"1001" when DATA_IN(17 downto 12)=b"100000" else
								b"1110" when DATA_IN(17 downto 12)=b"100010" else
								b"1111" when DATA_IN(17 downto 12)=b"100100" else
								b"0101" when DATA_IN(17 downto 12)=b"100110" else
								b"0010" when DATA_IN(17 downto 12)=b"101000" else
								b"1000" when DATA_IN(17 downto 12)=b"101010" else
								b"1100" when DATA_IN(17 downto 12)=b"101100" else
								b"0011" when DATA_IN(17 downto 12)=b"101110" else
								b"0111" when DATA_IN(17 downto 12)=b"110000" else
								b"0000" when DATA_IN(17 downto 12)=b"110010" else
								b"0100" when DATA_IN(17 downto 12)=b"110100" else
								b"1010" when DATA_IN(17 downto 12)=b"110110" else
								b"0001" when DATA_IN(17 downto 12)=b"111000" else
								b"1101" when DATA_IN(17 downto 12)=b"111010" else
								b"1011" when DATA_IN(17 downto 12)=b"111100" else
								b"0110" when DATA_IN(17 downto 12)=b"111110" else
								b"0100" when DATA_IN(17 downto 12)=b"100001" else
								b"0011" when DATA_IN(17 downto 12)=b"100011" else
								b"0010" when DATA_IN(17 downto 12)=b"100101" else
								b"1100" when DATA_IN(17 downto 12)=b"100111" else
								b"1001" when DATA_IN(17 downto 12)=b"101001" else
								b"0101" when DATA_IN(17 downto 12)=b"101011" else
								b"1111" when DATA_IN(17 downto 12)=b"101101" else
								b"1010" when DATA_IN(17 downto 12)=b"101111" else
								b"1011" when DATA_IN(17 downto 12)=b"110001" else
								b"1110" when DATA_IN(17 downto 12)=b"110011" else
								b"0001" when DATA_IN(17 downto 12)=b"110101" else
								b"0111" when DATA_IN(17 downto 12)=b"110111" else
								b"0110" when DATA_IN(17 downto 12)=b"111001" else
								b"0000" when DATA_IN(17 downto 12)=b"111011" else
								b"1000" when DATA_IN(17 downto 12)=b"111101" else
								b"1101" when DATA_IN(17 downto 12)=b"111111" else
								(others=>'0');
--siódmy sbox		
DATA_OUT(7 downto 4)<=  b"0100" when DATA_IN(11 downto 6)=b"000000" else
								b"1011" when DATA_IN(11 downto 6)=b"000010" else
								b"0010" when DATA_IN(11 downto 6)=b"000100" else
								b"1110" when DATA_IN(11 downto 6)=b"000110" else
								b"1111" when DATA_IN(11 downto 6)=b"001000" else
								b"0000" when DATA_IN(11 downto 6)=b"001010" else
								b"1000" when DATA_IN(11 downto 6)=b"001100" else
								b"1101" when DATA_IN(11 downto 6)=b"001110" else
								b"0011" when DATA_IN(11 downto 6)=b"010000" else
								b"1100" when DATA_IN(11 downto 6)=b"010010" else
								b"1001" when DATA_IN(11 downto 6)=b"010100" else
								b"0111" when DATA_IN(11 downto 6)=b"010110" else
								b"0101" when DATA_IN(11 downto 6)=b"011000" else
								b"1010" when DATA_IN(11 downto 6)=b"011010" else
								b"0110" when DATA_IN(11 downto 6)=b"011100" else
								b"0001" when DATA_IN(11 downto 6)=b"011110" else
								b"1101" when DATA_IN(11 downto 6)=b"000001" else
								b"0000" when DATA_IN(11 downto 6)=b"000011" else
								b"1011" when DATA_IN(11 downto 6)=b"000101" else
								b"0111" when DATA_IN(11 downto 6)=b"000111" else
								b"0100" when DATA_IN(11 downto 6)=b"001001" else
								b"1001" when DATA_IN(11 downto 6)=b"001011" else
								b"0001" when DATA_IN(11 downto 6)=b"001101" else
								b"1010" when DATA_IN(11 downto 6)=b"001111" else
								b"1110" when DATA_IN(11 downto 6)=b"010001" else
								b"0011" when DATA_IN(11 downto 6)=b"010011" else
								b"0101" when DATA_IN(11 downto 6)=b"010101" else
								b"1100" when DATA_IN(11 downto 6)=b"010111" else
								b"0010" when DATA_IN(11 downto 6)=b"011001" else
								b"1111" when DATA_IN(11 downto 6)=b"011011" else
								b"1000" when DATA_IN(11 downto 6)=b"011101" else
								b"0110" when DATA_IN(11 downto 6)=b"011111" else
								b"0001" when DATA_IN(11 downto 6)=b"100000" else
								b"0100" when DATA_IN(11 downto 6)=b"100010" else
								b"1011" when DATA_IN(11 downto 6)=b"100100" else
								b"1101" when DATA_IN(11 downto 6)=b"100110" else
								b"1100" when DATA_IN(11 downto 6)=b"101000" else
								b"0011" when DATA_IN(11 downto 6)=b"101010" else
								b"0111" when DATA_IN(11 downto 6)=b"101100" else
								b"1110" when DATA_IN(11 downto 6)=b"101110" else
								b"1010" when DATA_IN(11 downto 6)=b"110000" else
								b"1111" when DATA_IN(11 downto 6)=b"110010" else
								b"0110" when DATA_IN(11 downto 6)=b"110100" else
								b"1000" when DATA_IN(11 downto 6)=b"110110" else
								b"0000" when DATA_IN(11 downto 6)=b"111000" else
								b"0101" when DATA_IN(11 downto 6)=b"111010" else
								b"1001" when DATA_IN(11 downto 6)=b"111100" else
								b"0010" when DATA_IN(11 downto 6)=b"111110" else
								b"0110" when DATA_IN(11 downto 6)=b"100001" else
								b"1011" when DATA_IN(11 downto 6)=b"100011" else
								b"1101" when DATA_IN(11 downto 6)=b"100101" else
								b"1000" when DATA_IN(11 downto 6)=b"100111" else
								b"0001" when DATA_IN(11 downto 6)=b"101001" else
								b"0100" when DATA_IN(11 downto 6)=b"101011" else
								b"1010" when DATA_IN(11 downto 6)=b"101101" else
								b"0111" when DATA_IN(11 downto 6)=b"101111" else
								b"1001" when DATA_IN(11 downto 6)=b"110001" else
								b"0101" when DATA_IN(11 downto 6)=b"110011" else
								b"0000" when DATA_IN(11 downto 6)=b"110101" else
								b"1111" when DATA_IN(11 downto 6)=b"110111" else
								b"1110" when DATA_IN(11 downto 6)=b"111001" else
								b"0010" when DATA_IN(11 downto 6)=b"111011" else
								b"0011" when DATA_IN(11 downto 6)=b"111101" else
								b"1100" when DATA_IN(11 downto 6)=b"111111" else
								(others=>'0');
--ósmy sbox				
DATA_OUT(3 downto 0)<=  b"1101" when DATA_IN(5 downto 0)=b"000000" else
								b"0010" when DATA_IN(5 downto 0)=b"000010" else
								b"1000" when DATA_IN(5 downto 0)=b"000100" else
								b"0100" when DATA_IN(5 downto 0)=b"000110" else
								b"0110" when DATA_IN(5 downto 0)=b"001000" else
								b"1111" when DATA_IN(5 downto 0)=b"001010" else
								b"1011" when DATA_IN(5 downto 0)=b"001100" else
								b"0001" when DATA_IN(5 downto 0)=b"001110" else
								b"1010" when DATA_IN(5 downto 0)=b"010000" else
								b"1001" when DATA_IN(5 downto 0)=b"010010" else
								b"0011" when DATA_IN(5 downto 0)=b"010100" else
								b"1110" when DATA_IN(5 downto 0)=b"010110" else
								b"0101" when DATA_IN(5 downto 0)=b"011000" else
								b"0000" when DATA_IN(5 downto 0)=b"011010" else
								b"1100" when DATA_IN(5 downto 0)=b"011100" else
								b"0111" when DATA_IN(5 downto 0)=b"011110" else
								b"0001" when DATA_IN(5 downto 0)=b"000001" else
								b"1111" when DATA_IN(5 downto 0)=b"000011" else
								b"1101" when DATA_IN(5 downto 0)=b"000101" else
								b"1000" when DATA_IN(5 downto 0)=b"000111" else
								b"1010" when DATA_IN(5 downto 0)=b"001001" else
								b"0011" when DATA_IN(5 downto 0)=b"001011" else
								b"0111" when DATA_IN(5 downto 0)=b"001101" else
								b"0100" when DATA_IN(5 downto 0)=b"001111" else
								b"1100" when DATA_IN(5 downto 0)=b"010001" else
								b"0101" when DATA_IN(5 downto 0)=b"010011" else
								b"0110" when DATA_IN(5 downto 0)=b"010101" else
								b"1011" when DATA_IN(5 downto 0)=b"010111" else
								b"0000" when DATA_IN(5 downto 0)=b"011001" else
								b"1110" when DATA_IN(5 downto 0)=b"011011" else
								b"1001" when DATA_IN(5 downto 0)=b"011101" else
								b"0010" when DATA_IN(5 downto 0)=b"011111" else
								b"0111" when DATA_IN(5 downto 0)=b"100000" else
								b"1011" when DATA_IN(5 downto 0)=b"100010" else
								b"0100" when DATA_IN(5 downto 0)=b"100100" else
								b"0001" when DATA_IN(5 downto 0)=b"100110" else
								b"1001" when DATA_IN(5 downto 0)=b"101000" else
								b"1100" when DATA_IN(5 downto 0)=b"101010" else
								b"1110" when DATA_IN(5 downto 0)=b"101100" else
								b"0010" when DATA_IN(5 downto 0)=b"101110" else
								b"0000" when DATA_IN(5 downto 0)=b"110000" else
								b"0110" when DATA_IN(5 downto 0)=b"110010" else
								b"1010" when DATA_IN(5 downto 0)=b"110100" else
								b"1101" when DATA_IN(5 downto 0)=b"110110" else
								b"1111" when DATA_IN(5 downto 0)=b"111000" else
								b"1100" when DATA_IN(5 downto 0)=b"111010" else
								b"0101" when DATA_IN(5 downto 0)=b"111100" else
								b"1000" when DATA_IN(5 downto 0)=b"111110" else
								b"0010" when DATA_IN(5 downto 0)=b"100001" else
								b"0001" when DATA_IN(5 downto 0)=b"100011" else
								b"1110" when DATA_IN(5 downto 0)=b"100101" else
								b"0111" when DATA_IN(5 downto 0)=b"100111" else
								b"0100" when DATA_IN(5 downto 0)=b"101001" else
								b"1010" when DATA_IN(5 downto 0)=b"101011" else
								b"1000" when DATA_IN(5 downto 0)=b"101101" else
								b"1101" when DATA_IN(5 downto 0)=b"101111" else
								b"1111" when DATA_IN(5 downto 0)=b"110001" else
								b"1100" when DATA_IN(5 downto 0)=b"110011" else
								b"1001" when DATA_IN(5 downto 0)=b"110101" else
								b"0000" when DATA_IN(5 downto 0)=b"110111" else
								b"0011" when DATA_IN(5 downto 0)=b"111001" else
								b"0101" when DATA_IN(5 downto 0)=b"111011" else
								b"0110" when DATA_IN(5 downto 0)=b"111101" else
								b"1011" when DATA_IN(5 downto 0)=b"111111" else
								(others=>'0');
								
END ARCHITECTURE;