LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY LFSR IS PORT
(
CLK :IN STD_LOGIC;
INIT :IN STD_LOGIC;
DOUT :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END ENTITY;
ARCHITECTURE ARCH_LFSR OF LFSR IS
SIGNAL ISTATE : STD_LOGIC_VECTOR(63 DOWNTO 0);
BEGIN

PROCESS(CLK)
BEGIN
IF (INIT = '1') THEN ISTATE <= B"0000000000000000000000000000000000000000000000000000000000000001";
ELSIF(CLK'EVENT AND CLK = '1') THEN
--ISTATE <= ISTATE(62 DOWNTO 0) & (ISTATE(63) XOR ISTATE(3) XOR ISTATE(2) XOR ISTATE(0));
ISTATE(63 downto 1) <= ISTATE(62 DOWNTO 0) ;
ISTATE(0) <= (ISTATE(63) XOR ISTATE(3) XOR ISTATE(2) XOR ISTATE(0));
END IF;
END PROCESS;

DOUT <= ISTATE;
END ARCHITECTURE;