LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY PC_1 IS PORT
(
A :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
Y :OUT STD_LOGIC_VECTOR(55 DOWNTO 0)
);
END PC_1;
ARCHITECTURE ARCH_PC_1 OF PC_1 IS
BEGIN
Y(55)<=A(7);
Y(54)<=A(15);
Y(53)<=A(23);
Y(52)<=A(31);
Y(51)<=A(39);
Y(50)<=A(47);
Y(49)<=A(55);
Y(48)<=A(63);
Y(47)<=A(6);
Y(46)<=A(14);
Y(45)<=A(22);
Y(44)<=A(30);
Y(43)<=A(38);
Y(42)<=A(46);
Y(41)<=A(54);
Y(40)<=A(62);
Y(39)<=A(5);
Y(38)<=A(13);
Y(37)<=A(21);
Y(36)<=A(29);
Y(35)<=A(37);
Y(34)<=A(45);
Y(33)<=A(53);
Y(32)<=A(61);
Y(31)<=A(4);
Y(30)<=A(12);
Y(29)<=A(20);
Y(28)<=A(28);
Y(27)<=A(1);
Y(26)<=A(9);
Y(25)<=A(17);
Y(24)<=A(25);
Y(23)<=A(33);
Y(22)<=A(41);
Y(21)<=A(49);
Y(20)<=A(57);
Y(19)<=A(2);
Y(18)<=A(10);
Y(17)<=A(18);
Y(16)<=A(26);
Y(15)<=A(34);
Y(14)<=A(42);
Y(13)<=A(50);
Y(12)<=A(58);
Y(11)<=A(3);
Y(10)<=A(11);
Y(9)<=A(19);
Y(8)<=A(27);
Y(7)<=A(35);
Y(6)<=A(43);
Y(5)<=A(51);
Y(4)<=A(59);
Y(3)<=A(36);
Y(2)<=A(44);
Y(1)<=A(52);
Y(0)<=A(60);
END ARCHITECTURE;