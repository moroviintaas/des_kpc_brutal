LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY final_permutation IS PORT
(
A :IN STD_LOGIC_VECTOR(63 DOWNTO 0);
Y :OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
);
END final_permutation;
ARCHITECTURE ARCH_final_permutation OF final_permutation IS
BEGIN
Y(63)<=A(24);
Y(62)<=A(56);
Y(61)<=A(16);
Y(60)<=A(48);
Y(59)<=A(8);
Y(58)<=A(40);
Y(57)<=A(0);
Y(56)<=A(32);
Y(55)<=A(25);
Y(54)<=A(57);
Y(53)<=A(17);
Y(52)<=A(49);
Y(51)<=A(9);
Y(50)<=A(41);
Y(49)<=A(1);
Y(48)<=A(33);
Y(47)<=A(26);
Y(46)<=A(58);
Y(45)<=A(18);
Y(44)<=A(50);
Y(43)<=A(10);
Y(42)<=A(42);
Y(41)<=A(2);
Y(40)<=A(34);
Y(39)<=A(27);
Y(38)<=A(59);
Y(37)<=A(19);
Y(36)<=A(51);
Y(35)<=A(11);
Y(34)<=A(43);
Y(33)<=A(3);
Y(32)<=A(35);
Y(31)<=A(28);
Y(30)<=A(60);
Y(29)<=A(20);
Y(28)<=A(52);
Y(27)<=A(12);
Y(26)<=A(44);
Y(25)<=A(4);
Y(24)<=A(36);
Y(23)<=A(29);
Y(22)<=A(61);
Y(21)<=A(21);
Y(20)<=A(53);
Y(19)<=A(13);
Y(18)<=A(45);
Y(17)<=A(5);
Y(16)<=A(37);
Y(15)<=A(30);
Y(14)<=A(62);
Y(13)<=A(22);
Y(12)<=A(54);
Y(11)<=A(14);
Y(10)<=A(46);
Y(9)<=A(6);
Y(8)<=A(38);
Y(7)<=A(31);
Y(6)<=A(63);
Y(5)<=A(23);
Y(4)<=A(55);
Y(3)<=A(15);
Y(2)<=A(47);
Y(1)<=A(7);
Y(0)<=A(39);
END ARCHITECTURE;